*** SPICE deck for cell 2bit_multiplier2{lay} from library ServetCelik_ELE419_Project
*** Created on Sal Oca 02, 2024 01:28:45
*** Last revised on Cmt Oca 13, 2024 16:23:06
*** Written on Cmt Oca 13, 2024 16:23:09 by Electric VLSI Design System, version 9.07
*** Layout tech: mocmos, foundry MOSIS
*** UC SPICE *** , MIN_RESIST 4.0, MIN_CAPAC 0.1FF

*** SUBCIRCUIT ServetCelik_ELE419_Project__NAND_gate2 FROM CELL NAND_gate2{lay}
.SUBCKT ServetCelik_ELE419_Project__NAND_gate2 0 A A_nand_B B vdd
Mnmos_0 net_34 B A_nand_B 0 N L=0.6U W=2.4U AS=4.56P AD=1.418P PS=7.3U PD=4.05U
Mnmos_1 0 A net_34 0 N L=0.6U W=2.4U AS=1.418P AD=16.83P PS=4.05U PD=27.9U
Mpmos_0 A_nand_B A vdd vdd P L=0.6U W=2.4U AS=13.05P AD=4.56P PS=21U PD=7.3U
Mpmos_1 vdd B A_nand_B vdd P L=0.6U W=2.4U AS=4.56P AD=13.05P PS=7.3U PD=21U
.ENDS ServetCelik_ELE419_Project__NAND_gate2

*** SUBCIRCUIT ServetCelik_ELE419_Project__inverter2 FROM CELL inverter2{lay}
.SUBCKT ServetCelik_ELE419_Project__inverter2 0 A A_not vdd
Mnmos_0 A_not A 0 0 N L=0.6U W=1.2U AS=9.54P AD=4.725P PS=18.9U PD=9U
Mpmos_0 A_not A vdd vdd P L=0.6U W=2.4U AS=12.33P AD=4.725P PS=21.9U PD=9U
.ENDS ServetCelik_ELE419_Project__inverter2

*** SUBCIRCUIT ServetCelik_ELE419_Project__AND_gate2 FROM CELL AND_gate2{lay}
.SUBCKT ServetCelik_ELE419_Project__AND_gate2 0 A A_and_B B vdd
XNAND_gat_2 0 A net_0 B vdd ServetCelik_ELE419_Project__NAND_gate2
Xinverter_2 0 net_0 A_and_B vdd ServetCelik_ELE419_Project__inverter2
.ENDS ServetCelik_ELE419_Project__AND_gate2

*** SUBCIRCUIT ServetCelik_ELE419_Project__XOR_gate2 FROM CELL XOR_gate2{lay}
.SUBCKT ServetCelik_ELE419_Project__XOR_gate2 0 A A_xor_B B vdd
Mnmos_7 net_258 B 0 0 N L=0.6U W=1.2U AS=5.783P AD=1.845P PS=11.7U PD=4.2U
Mnmos_8 A_xor_B A net_258 0 N L=0.6U W=1.2U AS=1.845P AD=2.858P PS=4.2U PD=5.1U
Mnmos_9 net_259 net_263 A_xor_B 0 N L=0.6U W=1.2U AS=2.858P AD=2.025P PS=5.1U PD=4.5U
Mnmos_10 0 net_230 net_259 0 N L=0.6U W=1.2U AS=2.025P AD=5.783P PS=4.5U PD=11.7U
Mnmos_11 net_263 A 0 0 N L=0.6U W=1.2U AS=5.783P AD=4.185P PS=11.7U PD=8.4U
Mnmos_12 net_230 B 0 0 N L=0.6U W=1.2U AS=5.783P AD=4.725P PS=11.7U PD=9U
Mpmos_10 A_xor_B B net_199 vdd P L=0.6U W=2.4U AS=4.995P AD=2.858P PS=8.1U PD=5.1U
Mpmos_11 net_199 A A_xor_B vdd P L=0.6U W=2.4U AS=2.858P AD=4.995P PS=5.1U PD=8.1U
Mpmos_12 vdd net_263 net_199 vdd P L=0.6U W=2.4U AS=4.995P AD=7.808P PS=8.1U PD=12.6U
Mpmos_13 net_199 net_230 vdd vdd P L=0.6U W=2.4U AS=7.808P AD=4.995P PS=12.6U PD=8.1U
Mpmos_14 net_263 A vdd vdd P L=0.6U W=2.4U AS=7.808P AD=4.185P PS=12.6U PD=8.4U
Mpmos_15 net_230 B vdd vdd P L=0.6U W=2.4U AS=7.808P AD=4.725P PS=12.6U PD=9U
.ENDS ServetCelik_ELE419_Project__XOR_gate2

*** SUBCIRCUIT ServetCelik_ELE419_Project__halfAdder2 FROM CELL halfAdder2{lay}
.SUBCKT ServetCelik_ELE419_Project__halfAdder2 0 A B halfAdder_carry halfAdder_sum vdd
XAND_gate_2 0 A halfAdder_carry B vdd ServetCelik_ELE419_Project__AND_gate2
XXOR_gate_2 0 A halfAdder_sum B vdd ServetCelik_ELE419_Project__XOR_gate2
.ENDS ServetCelik_ELE419_Project__halfAdder2

*** TOP LEVEL CELL: 2bit_multiplier2{lay}
XAND_gate_4 0 A1 net_18 B1 vdd ServetCelik_ELE419_Project__AND_gate2
XAND_gate_5 0 A0 net_11 B1 vdd ServetCelik_ELE419_Project__AND_gate2
XAND_gate_6 0 A1 net_0 B0 vdd ServetCelik_ELE419_Project__AND_gate2
XAND_gate_7 0 A0 P0 B0 vdd ServetCelik_ELE419_Project__AND_gate2
XhalfAdde_2 0 net_11 net_0 net_21 P1 vdd ServetCelik_ELE419_Project__halfAdder2
XhalfAdde_3 0 net_18 net_21 P3 P2 vdd ServetCelik_ELE419_Project__halfAdder2

* Spice Code nodes in cell cell '2bit_multiplier2{lay}'
vdd vdd 0 DC 5
VinA1 A1 0 DC 0
VinA0 A0 0 DC 0
VinB1 B1 0 DC 5
VinB0 B0 0 DC 5
.tran 10u 40u
* Trailer cards are described in this file:
.INC C:\Users\Servet\Desktop\C5_models.txt
.END
