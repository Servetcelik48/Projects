*** SPICE deck for cell Analog_barepadframe_1.5mmX1.5mm{lay} from library ServetCelik_ELE419_Project
*** Created on Çar May 27, 2009 02:00:56
*** Last revised on Sal Oca 16, 2024 13:00:02
*** Written on Sal Oca 16, 2024 13:01:42 by Electric VLSI Design System, version 9.07
*** Layout tech: mocmos, foundry MOSIS
*** UC SPICE *** , MIN_RESIST 4.0, MIN_CAPAC 0.1FF

*** SUBCIRCUIT ServetCelik_ELE419_Project__NOR_gate2 FROM CELL NOR_gate2{lay}
.SUBCKT ServetCelik_ELE419_Project__NOR_gate2 0 A A_nor_B B vdd
Mnmos_2 A_nor_B A 0 0 N L=0.6U W=1.2U AS=6.525P AD=3.21P PS=13.5U PD=6.1U
Mnmos_3 0 B A_nor_B 0 N L=0.6U W=1.2U AS=3.21P AD=6.525P PS=6.1U PD=13.5U
Mpmos_2 net_75 A vdd vdd P L=0.6U W=2.4U AS=13.05P AD=1.418P PS=22.5U PD=4.05U
Mpmos_3 A_nor_B B net_75 vdd P L=0.6U W=2.4U AS=1.418P AD=3.21P PS=4.05U PD=6.1U
.ENDS ServetCelik_ELE419_Project__NOR_gate2

*** SUBCIRCUIT ServetCelik_ELE419_Project__inverter2 FROM CELL inverter2{lay}
.SUBCKT ServetCelik_ELE419_Project__inverter2 0 A A_not vdd
Mnmos_0 A_not A 0 0 N L=0.6U W=1.2U AS=9.54P AD=4.725P PS=18.9U PD=9U
Mpmos_0 A_not A vdd vdd P L=0.6U W=2.4U AS=12.33P AD=4.725P PS=21.9U PD=9U
.ENDS ServetCelik_ELE419_Project__inverter2

*** SUBCIRCUIT ServetCelik_ELE419_Project__OR_gate2 FROM CELL OR_gate2{lay}
.SUBCKT ServetCelik_ELE419_Project__OR_gate2 0 A A_or_B B vdd
XNOR_gate_2 0 A net_30 B vdd ServetCelik_ELE419_Project__NOR_gate2
Xinverter_1 0 net_30 A_or_B vdd ServetCelik_ELE419_Project__inverter2
.ENDS ServetCelik_ELE419_Project__OR_gate2

*** SUBCIRCUIT ServetCelik_ELE419_Project__NAND_gate2 FROM CELL NAND_gate2{lay}
.SUBCKT ServetCelik_ELE419_Project__NAND_gate2 0 A A_nand_B B vdd
Mnmos_0 net_34 B A_nand_B 0 N L=0.6U W=2.4U AS=4.56P AD=1.418P PS=7.3U PD=4.05U
Mnmos_1 0 A net_34 0 N L=0.6U W=2.4U AS=1.418P AD=16.83P PS=4.05U PD=27.9U
Mpmos_0 A_nand_B A vdd vdd P L=0.6U W=2.4U AS=13.05P AD=4.56P PS=21U PD=7.3U
Mpmos_1 vdd B A_nand_B vdd P L=0.6U W=2.4U AS=4.56P AD=13.05P PS=7.3U PD=21U
.ENDS ServetCelik_ELE419_Project__NAND_gate2

*** SUBCIRCUIT ServetCelik_ELE419_Project__AND_gate2 FROM CELL AND_gate2{lay}
.SUBCKT ServetCelik_ELE419_Project__AND_gate2 0 A A_and_B B vdd
XNAND_gat_2 0 A net_0 B vdd ServetCelik_ELE419_Project__NAND_gate2
Xinverter_2 0 net_0 A_and_B vdd ServetCelik_ELE419_Project__inverter2
.ENDS ServetCelik_ELE419_Project__AND_gate2

*** SUBCIRCUIT ServetCelik_ELE419_Project__XOR_gate2 FROM CELL XOR_gate2{lay}
.SUBCKT ServetCelik_ELE419_Project__XOR_gate2 0 A A_xor_B B vdd
Mnmos_7 net_258 B 0 0 N L=0.6U W=1.2U AS=5.783P AD=1.845P PS=11.7U PD=4.2U
Mnmos_8 A_xor_B A net_258 0 N L=0.6U W=1.2U AS=1.845P AD=2.858P PS=4.2U PD=5.1U
Mnmos_9 net_259 net_263 A_xor_B 0 N L=0.6U W=1.2U AS=2.858P AD=2.025P PS=5.1U PD=4.5U
Mnmos_10 0 net_230 net_259 0 N L=0.6U W=1.2U AS=2.025P AD=5.783P PS=4.5U PD=11.7U
Mnmos_11 net_263 A 0 0 N L=0.6U W=1.2U AS=5.783P AD=4.185P PS=11.7U PD=8.4U
Mnmos_12 net_230 B 0 0 N L=0.6U W=1.2U AS=5.783P AD=4.725P PS=11.7U PD=9U
Mpmos_10 A_xor_B B net_199 vdd P L=0.6U W=2.4U AS=4.995P AD=2.858P PS=8.1U PD=5.1U
Mpmos_11 net_199 A A_xor_B vdd P L=0.6U W=2.4U AS=2.858P AD=4.995P PS=5.1U PD=8.1U
Mpmos_12 vdd net_263 net_199 vdd P L=0.6U W=2.4U AS=4.995P AD=7.808P PS=8.1U PD=12.6U
Mpmos_13 net_199 net_230 vdd vdd P L=0.6U W=2.4U AS=7.808P AD=4.995P PS=12.6U PD=8.1U
Mpmos_14 net_263 A vdd vdd P L=0.6U W=2.4U AS=7.808P AD=4.185P PS=12.6U PD=8.4U
Mpmos_15 net_230 B vdd vdd P L=0.6U W=2.4U AS=7.808P AD=4.725P PS=12.6U PD=9U
.ENDS ServetCelik_ELE419_Project__XOR_gate2

*** SUBCIRCUIT ServetCelik_ELE419_Project__halfAdder2 FROM CELL halfAdder2{lay}
.SUBCKT ServetCelik_ELE419_Project__halfAdder2 0 A B halfAdder_carry halfAdder_sum vdd
XAND_gate_2 0 A halfAdder_carry B vdd ServetCelik_ELE419_Project__AND_gate2
XXOR_gate_2 0 A halfAdder_sum B vdd ServetCelik_ELE419_Project__XOR_gate2
.ENDS ServetCelik_ELE419_Project__halfAdder2

*** SUBCIRCUIT ServetCelik_ELE419_Project__fullAdder2 FROM CELL fullAdder2{lay}
.SUBCKT ServetCelik_ELE419_Project__fullAdder2 0 A B Cin fullAdder_carry fullAdder_sum vdd
XOR_gate2_0 0 net_39 fullAdder_carry net_42 vdd ServetCelik_ELE419_Project__OR_gate2
XhalfAdde_2 0 net_47 Cin net_42 fullAdder_sum vdd ServetCelik_ELE419_Project__halfAdder2
XhalfAdde_3 0 A B net_39 net_47 vdd ServetCelik_ELE419_Project__halfAdder2
.ENDS ServetCelik_ELE419_Project__fullAdder2

*** SUBCIRCUIT ServetCelik_ELE419_Project__2bit_RCA2 FROM CELL 2bit_RCA2{lay}
.SUBCKT ServetCelik_ELE419_Project__2bit_RCA2 0 A0 A1 B0 B1 carry S0 S1 vdd
XfullAdde_2 0 A1 B1 net_34 carry S1 vdd ServetCelik_ELE419_Project__fullAdder2
XfullAdde_3 0 A0 B0 0 net_34 S0 vdd ServetCelik_ELE419_Project__fullAdder2
.ENDS ServetCelik_ELE419_Project__2bit_RCA2

*** SUBCIRCUIT ServetCelik_ELE419_Project__2bit_multiplier2 FROM CELL 2bit_multiplier2{lay}
.SUBCKT ServetCelik_ELE419_Project__2bit_multiplier2 0 A0 A1 B0 B1 P0 P1 P2 P3 vdd
XAND_gate_4 0 A1 net_18 B1 vdd ServetCelik_ELE419_Project__AND_gate2
XAND_gate_5 0 A0 net_11 B1 vdd ServetCelik_ELE419_Project__AND_gate2
XAND_gate_6 0 A1 net_0 B0 vdd ServetCelik_ELE419_Project__AND_gate2
XAND_gate_7 0 A0 P0 B0 vdd ServetCelik_ELE419_Project__AND_gate2
XhalfAdde_2 0 net_11 net_0 net_21 P1 vdd ServetCelik_ELE419_Project__halfAdder2
XhalfAdde_3 0 net_18 net_21 P3 P2 vdd ServetCelik_ELE419_Project__halfAdder2
.ENDS ServetCelik_ELE419_Project__2bit_multiplier2

*** SUBCIRCUIT ServetCelik_ELE419_Project__4bit_RCA2 FROM CELL 4bit_RCA2{lay}
.SUBCKT ServetCelik_ELE419_Project__4bit_RCA2 0 A0 A1 A2 A3 B0 B1 B2 B3 carry S0 S1 S2 S3 vdd
XfullAdde_4 0 A1 B1 net_175 net_106 S1 vdd ServetCelik_ELE419_Project__fullAdder2
XfullAdde_5 0 A0 B0 0 net_175 S0 vdd ServetCelik_ELE419_Project__fullAdder2
XfullAdde_8 0 A3 B3 net_208 carry S3 vdd ServetCelik_ELE419_Project__fullAdder2
XfullAdde_9 0 A2 B2 net_106 net_208 S2 vdd ServetCelik_ELE419_Project__fullAdder2
.ENDS ServetCelik_ELE419_Project__4bit_RCA2

*** SUBCIRCUIT ServetCelik_ELE419_Project__4bit_multiplier2 FROM CELL 4bit_multiplier2{lay}
.SUBCKT ServetCelik_ELE419_Project__4bit_multiplier2 0 A0 A1 A2 A3 B0 B1 B2 B3 carry P0 P1 P2 P3 P4 P5 P6 P7 vdd
X2bit_RCA_1 0 net_762 net_755 net_771 net_783 carry P6 P7 vdd ServetCelik_ELE419_Project__2bit_RCA2
X2bit_mul_4 0 A2 A3 B2 B3 net_369 net_364 net_771 net_783 vdd ServetCelik_ELE419_Project__2bit_multiplier2
X2bit_mul_5 0 A0 A1 B2 B3 net_249 net_258 net_311 net_316 vdd ServetCelik_ELE419_Project__2bit_multiplier2
X2bit_mul_6 0 A2 A3 B0 B1 net_288 net_291 net_296 net_299 vdd ServetCelik_ELE419_Project__2bit_multiplier2
X2bit_mul_7 0 A0 A1 B0 B1 P0 P1 net_350 net_353 vdd ServetCelik_ELE419_Project__2bit_multiplier2
X4bit_RCA_2 0 net_288 net_291 net_296 net_299 net_249 net_258 net_311 net_316 net_752 net_322 net_326 net_330 net_335 vdd ServetCelik_ELE419_Project__4bit_RCA2
X4bit_RCA_3 0 net_350 net_353 net_369 net_364 net_322 net_326 net_330 net_335 net_743 P2 P3 P4 P5 vdd ServetCelik_ELE419_Project__4bit_RCA2
XhalfAdde_2 0 net_752 net_743 net_755 net_762 vdd ServetCelik_ELE419_Project__halfAdder2
.ENDS ServetCelik_ELE419_Project__4bit_multiplier2

*** SUBCIRCUIT ServetCelik_ELE419_Project__8bit_RCA2 FROM CELL 8bit_RCA2{lay}
.SUBCKT ServetCelik_ELE419_Project__8bit_RCA2 0 A0 A1 A2 A3 A4 A5 A6 A7 B0 B1 B2 B3 B4 B5 B6 B7 carry S0 S1 S2 S3 S4 S5 S6 S7 vdd
XfullAdde_8 0 A1 B1 net_139 net_126 S1 vdd ServetCelik_ELE419_Project__fullAdder2
XfullAdde_9 0 A0 B0 0 net_139 S0 vdd ServetCelik_ELE419_Project__fullAdder2
XfullAdde_10 0 A3 B3 net_165 net_263 S3 vdd ServetCelik_ELE419_Project__fullAdder2
XfullAdde_11 0 A2 B2 net_126 net_165 S2 vdd ServetCelik_ELE419_Project__fullAdder2
XfullAdde_12 0 A5 B5 net_209 net_196 S5 vdd ServetCelik_ELE419_Project__fullAdder2
XfullAdde_13 0 A4 B4 net_263 net_209 S4 vdd ServetCelik_ELE419_Project__fullAdder2
XfullAdde_14 0 A7 B7 net_235 carry S7 vdd ServetCelik_ELE419_Project__fullAdder2
XfullAdde_15 0 A6 B6 net_196 net_235 S6 vdd ServetCelik_ELE419_Project__fullAdder2
.ENDS ServetCelik_ELE419_Project__8bit_RCA2

*** SUBCIRCUIT ServetCelik_ELE419_Project__8bit_multiplier2 FROM CELL 8bit_multiplier2{lay}
.SUBCKT ServetCelik_ELE419_Project__8bit_multiplier2 0 A0 A1 A2 A3 A4 A5 A6 A7 B0 B1 B2 B3 B4 B5 B6 B7 P0 P1 P10 P11 P12 P13 P14 P15 P2 P3 P4 P5 P6 P7 P8 P9 vdd
X4bit_mul_4 0 A4 A5 A6 A7 B0 B1 B2 B3 4bit_mul_4_carry net_77 net_81 net_82 net_83 net_84 net_85 net_101 net_105 vdd ServetCelik_ELE419_Project__4bit_multiplier2
X4bit_mul_5 0 A4 A5 A6 A7 B4 B5 B6 B7 4bit_mul_5_carry net_257 net_264 net_273 net_277 net_281 net_285 net_292 net_718 vdd ServetCelik_ELE419_Project__4bit_multiplier2
X4bit_mul_6 0 A0 A1 A2 A3 B0 B1 B2 B3 4bit_mul_6_carry P0 P1 P2 P3 net_111 net_119 net_116 net_122 vdd ServetCelik_ELE419_Project__4bit_multiplier2
X4bit_mul_7 0 A0 A1 A2 A3 B4 B5 B6 B7 4bit_mul_7_carry net_7 net_4 net_15 net_18 net_22 net_26 net_30 net_33 vdd ServetCelik_ELE419_Project__4bit_multiplier2
X8bit_RCA_3 0 net_237 net_240 net_245 net_246 net_255 0 0 0 net_257 net_264 net_273 net_277 net_281 net_285 net_292 net_718 8bit_RCA_3_carry P8 P9 P10 P11 P12 P13 P14 P15 vdd ServetCelik_ELE419_Project__8bit_RCA2
X8bit_RCA_4 0 net_7 net_4 net_15 net_18 net_22 net_26 net_30 net_33 net_77 net_81 net_82 net_83 net_84 net_85 net_101 net_105 net_255 net_142 net_143 net_147 net_150 net_153 net_156 net_159 net_162 vdd ServetCelik_ELE419_Project__8bit_RCA2
X8bit_RCA_5 0 net_111 net_119 net_116 net_122 0 net_156 0 0 net_142 net_143 net_147 net_150 net_153 0 net_159 net_162 8bit_RCA_5_carry P4 P5 P6 P7 net_237 net_240 net_245 net_246 vdd ServetCelik_ELE419_Project__8bit_RCA2
.ENDS ServetCelik_ELE419_Project__8bit_multiplier2

*** SUBCIRCUIT MOSIS_SUBM_PADS_C5__Frame_Corner FROM CELL MOSIS_SUBM_PADS_C5:Frame_Corner{lay}
.SUBCKT MOSIS_SUBM_PADS_C5__Frame_Corner 0 gnd

* Spice Code nodes in cell cell 'MOSIS_SUBM_PADS_C5:Frame_Corner{lay}'
R1 vdd gnd 100G
.ENDS MOSIS_SUBM_PADS_C5__Frame_Corner

*** SUBCIRCUIT MOSIS_SUBM_PADS_C5__Nact_PWell_diode FROM CELL MOSIS_SUBM_PADS_C5:Nact_PWell_diode{lay}
.SUBCKT MOSIS_SUBM_PADS_C5__Nact_PWell_diode N_act P_well

* Spice Code nodes in cell cell 'MOSIS_SUBM_PADS_C5:Nact_PWell_diode{lay}'
D1 P_well N_act Dnpn
.model Dnpn D is=1e-18 n=1
.ENDS MOSIS_SUBM_PADS_C5__Nact_PWell_diode

*** SUBCIRCUIT MOSIS_SUBM_PADS_C5__Pact_Nwell_diode FROM CELL MOSIS_SUBM_PADS_C5:Pact_Nwell_diode{lay}
.SUBCKT MOSIS_SUBM_PADS_C5__Pact_Nwell_diode N_well P_act

* Spice Code nodes in cell cell 'MOSIS_SUBM_PADS_C5:Pact_Nwell_diode{lay}'
D2 P_act N_well Dpnp
.model Dpnp D is=1e-18 n=1
.ENDS MOSIS_SUBM_PADS_C5__Pact_Nwell_diode

*** SUBCIRCUIT MOSIS_SUBM_PADS_C5__Vdd_Gnd_bus FROM CELL MOSIS_SUBM_PADS_C5:Vdd_Gnd_bus{lay}
.SUBCKT MOSIS_SUBM_PADS_C5__Vdd_Gnd_bus 0 vdd_1

* Spice Code nodes in cell cell 'MOSIS_SUBM_PADS_C5:Vdd_Gnd_bus{lay}'
R1 vdd_1 gnd_1 10g
.ENDS MOSIS_SUBM_PADS_C5__Vdd_Gnd_bus

*** SUBCIRCUIT MOSIS_SUBM_PADS_C5__Pad_Analog FROM CELL MOSIS_SUBM_PADS_C5:Pad_Analog{lay}
.SUBCKT MOSIS_SUBM_PADS_C5__Pad_Analog 0 Analog vdd_1
XNact_PWe_0 Analog 0 MOSIS_SUBM_PADS_C5__Nact_PWell_diode
XNwell_Pa_0 vdd_1 Analog MOSIS_SUBM_PADS_C5__Pact_Nwell_diode
XVdd_Gnd__0 0 vdd_1 MOSIS_SUBM_PADS_C5__Vdd_Gnd_bus
.ENDS MOSIS_SUBM_PADS_C5__Pad_Analog

*** SUBCIRCUIT MOSIS_SUBM_PADS_C5__Pad_Gnd FROM CELL MOSIS_SUBM_PADS_C5:Pad_Gnd{lay}
.SUBCKT MOSIS_SUBM_PADS_C5__Pad_Gnd 0 dvdd
XBus_Vdd__0 0 dvdd MOSIS_SUBM_PADS_C5__Vdd_Gnd_bus
XNact_PWe_0 0 0 MOSIS_SUBM_PADS_C5__Nact_PWell_diode
XNwell_Pa_0 dvdd 0 MOSIS_SUBM_PADS_C5__Pact_Nwell_diode
.ENDS MOSIS_SUBM_PADS_C5__Pad_Gnd

*** SUBCIRCUIT MOSIS_SUBM_PADS_C5__Pad_Vdd FROM CELL MOSIS_SUBM_PADS_C5:Pad_Vdd{lay}
.SUBCKT MOSIS_SUBM_PADS_C5__Pad_Vdd 0 VDD_PAD
XBus_Vdd__1 0 VDD_PAD MOSIS_SUBM_PADS_C5__Vdd_Gnd_bus
XNact_PWe_0 VDD_PAD 0 MOSIS_SUBM_PADS_C5__Nact_PWell_diode
XNwell_Pa_0 VDD_PAD VDD_PAD MOSIS_SUBM_PADS_C5__Pact_Nwell_diode
.ENDS MOSIS_SUBM_PADS_C5__Pad_Vdd

*** TOP LEVEL CELL: Analog_barepadframe_1.5mmX1.5mm{lay}
X8bit_mul_0 8bit_mul_0_gnd 8bit_mul_0_A0 8bit_mul_0_A1 8bit_mul_0_A2 8bit_mul_0_A3 8bit_mul_0_A4 8bit_mul_0_A5 8bit_mul_0_A6 8bit_mul_0_A7 8bit_mul_0_B0 8bit_mul_0_B1 8bit_mul_0_B2 8bit_mul_0_B3 8bit_mul_0_B4 8bit_mul_0_B5 8bit_mul_0_B6 8bit_mul_0_B7 8bit_mul_0_P0 8bit_mul_0_P1 8bit_mul_0_P10 8bit_mul_0_P11 8bit_mul_0_P12 8bit_mul_0_P13 8bit_mul_0_P14 8bit_mul_0_P15 8bit_mul_0_P2 8bit_mul_0_P3 8bit_mul_0_P4 8bit_mul_0_P5 8bit_mul_0_P6 8bit_mul_0_P7 8bit_mul_0_P8 8bit_mul_0_P9 vdd 
+ServetCelik_ELE419_Project__8bit_multiplier2
XI_O_Corn_0 vdd 0 MOSIS_SUBM_PADS_C5__Frame_Corner
XI_O_Corn_1 vdd 0 MOSIS_SUBM_PADS_C5__Frame_Corner
XI_O_Corn_2 vdd 0 MOSIS_SUBM_PADS_C5__Frame_Corner
XI_O_Corn_3 vdd 0 MOSIS_SUBM_PADS_C5__Frame_Corner
XPAD_M3M2_17 0 Pin35 vdd MOSIS_SUBM_PADS_C5__Pad_Analog
XPAD_M3M2_18 0 Pin34 vdd MOSIS_SUBM_PADS_C5__Pad_Analog
XPAD_M3M2_19 0 Pin33 vdd MOSIS_SUBM_PADS_C5__Pad_Analog
XPAD_M3M2_20 0 Pin32 vdd MOSIS_SUBM_PADS_C5__Pad_Analog
XPAD_M3M2_21 0 Pin31 vdd MOSIS_SUBM_PADS_C5__Pad_Analog
XPAD_M3M2_22 0 Pin30 vdd MOSIS_SUBM_PADS_C5__Pad_Analog
XPAD_M3M2_23 0 Pin29 vdd MOSIS_SUBM_PADS_C5__Pad_Analog
XPAD_M3M2_24 0 Pin28 vdd MOSIS_SUBM_PADS_C5__Pad_Analog
XPAD_M3M2_25 0 Pin27 vdd MOSIS_SUBM_PADS_C5__Pad_Analog
XPAD_M3M2_26 0 Pin26 vdd MOSIS_SUBM_PADS_C5__Pad_Analog
XPAD_M3M2_45 0 Pin25 vdd MOSIS_SUBM_PADS_C5__Pad_Analog
XPAD_M3M2_60 0 Pin24 vdd MOSIS_SUBM_PADS_C5__Pad_Analog
XPAD_M3M2_75 0 Pin23 vdd MOSIS_SUBM_PADS_C5__Pad_Analog
XPAD_M3M2_90 0 Pin22 vdd MOSIS_SUBM_PADS_C5__Pad_Analog
XPAD_M3M2_105 0 Pin21 vdd MOSIS_SUBM_PADS_C5__Pad_Analog
XPAD_M3M2_135 0 Pin19 vdd MOSIS_SUBM_PADS_C5__Pad_Analog
XPAD_M3M2_150 0 Pin18 vdd MOSIS_SUBM_PADS_C5__Pad_Analog
XPAD_M3M2_165 0 Pin17 vdd MOSIS_SUBM_PADS_C5__Pad_Analog
XPAD_M3M2_180 0 Pin16 vdd MOSIS_SUBM_PADS_C5__Pad_Analog
XPAD_M3M2_212 0 Pin15 vdd MOSIS_SUBM_PADS_C5__Pad_Analog
XPAD_M3M2_213 0 Pin14 vdd MOSIS_SUBM_PADS_C5__Pad_Analog
XPAD_M3M2_214 0 Pin13 vdd MOSIS_SUBM_PADS_C5__Pad_Analog
XPAD_M3M2_215 0 Pin12 vdd MOSIS_SUBM_PADS_C5__Pad_Analog
XPAD_M3M2_216 0 Pin11 vdd MOSIS_SUBM_PADS_C5__Pad_Analog
XPAD_M3M2_217 0 Pin10 vdd MOSIS_SUBM_PADS_C5__Pad_Analog
XPAD_M3M2_218 0 Pin9 vdd MOSIS_SUBM_PADS_C5__Pad_Analog
XPAD_M3M2_219 0 Pin8 vdd MOSIS_SUBM_PADS_C5__Pad_Analog
XPAD_M3M2_220 0 Pin7 vdd MOSIS_SUBM_PADS_C5__Pad_Analog
XPAD_M3M2_221 0 Pin6 vdd MOSIS_SUBM_PADS_C5__Pad_Analog
XPAD_M3M2_222 0 AAAAA vdd MOSIS_SUBM_PADS_C5__Pad_Analog
XPAD_M3M2_224 0 Pin39 vdd MOSIS_SUBM_PADS_C5__Pad_Analog
XPAD_M3M2_225 0 Pin38 vdd MOSIS_SUBM_PADS_C5__Pad_Analog
XPAD_M3M2_226 0 Pin37 vdd MOSIS_SUBM_PADS_C5__Pad_Analog
XPAD_M3M2_227 0 Pin36 vdd MOSIS_SUBM_PADS_C5__Pad_Analog
XPAD_M3M2_228 0 Pin5 vdd MOSIS_SUBM_PADS_C5__Pad_Analog
XPAD_M3M2_229 0 Pin4 vdd MOSIS_SUBM_PADS_C5__Pad_Analog
XPAD_M3M2_230 0 Pin3 vdd MOSIS_SUBM_PADS_C5__Pad_Analog
XPAD_M3M2_231 0 Pin2 vdd MOSIS_SUBM_PADS_C5__Pad_Analog
XPad_Gnd_0 0 vdd MOSIS_SUBM_PADS_C5__Pad_Gnd
XPad_Vdd_0 0 vdd MOSIS_SUBM_PADS_C5__Pad_Vdd

* Spice Code nodes in cell cell 'Analog_barepadframe_1.5mmX1.5mm{lay}'
vdd vdd 0 DC 5
VinPin1 Pin1 0 DC 5
VinA6 A6 0 DC 5
VinA5 A5 0 DC 5
VinA4 A4 0 DC 5
VinA3 A3 0 DC 5
VinA2 A2 0 DC 5
VinA1 A1 0 DC 5
VinA0 A0 0 DC 5
VinB7 B7 0 DC 5
VinB6 B6 0 DC 5
VinB5 B5 0 DC 0
VinB4 B4 0 DC 5
VinB3 B3 0 DC 5
VinB2 B2 0 DC 5
VinB1 B1 0 DC 0
VinB0 B0 0 DC 5
.tran 10u 40u
* Trailer cards are described in this file:
.INC C:\Users\Servet\Desktop\C5_models.txt
.END
