*** SPICE deck for cell 8bit_ALU{lay} from library ServetCelik_ELE419_Project
*** Created on Pzt Oca 15, 2024 12:52:19
*** Last revised on Çar Oca 17, 2024 18:08:42
*** Written on Per Oca 18, 2024 09:23:30 by Electric VLSI Design System, version 9.07
*** Layout tech: mocmos, foundry MOSIS
*** UC SPICE *** , MIN_RESIST 4.0, MIN_CAPAC 0.1FF

*** SUBCIRCUIT ServetCelik_ELE419_Project__NOR_gate2 FROM CELL NOR_gate2{lay}
.SUBCKT ServetCelik_ELE419_Project__NOR_gate2 0 A A_nor_B B vdd
Mnmos_2 A_nor_B A 0 0 N L=0.6U W=1.2U AS=6.525P AD=3.21P PS=13.5U PD=6.1U
Mnmos_3 0 B A_nor_B 0 N L=0.6U W=1.2U AS=3.21P AD=6.525P PS=6.1U PD=13.5U
Mpmos_2 net_75 A vdd vdd P L=0.6U W=2.4U AS=13.05P AD=1.418P PS=22.5U PD=4.05U
Mpmos_3 A_nor_B B net_75 vdd P L=0.6U W=2.4U AS=1.418P AD=3.21P PS=4.05U PD=6.1U
.ENDS ServetCelik_ELE419_Project__NOR_gate2

*** SUBCIRCUIT ServetCelik_ELE419_Project__inverter2 FROM CELL inverter2{lay}
.SUBCKT ServetCelik_ELE419_Project__inverter2 0 A A_not vdd
Mnmos_0 A_not A 0 0 N L=0.6U W=1.2U AS=9.54P AD=4.725P PS=18.9U PD=9U
Mpmos_0 A_not A vdd vdd P L=0.6U W=2.4U AS=12.33P AD=4.725P PS=21.9U PD=9U
.ENDS ServetCelik_ELE419_Project__inverter2

*** SUBCIRCUIT ServetCelik_ELE419_Project__OR_gate2 FROM CELL OR_gate2{lay}
.SUBCKT ServetCelik_ELE419_Project__OR_gate2 0 A A_or_B B vdd
XNOR_gate_2 0 A net_30 B vdd ServetCelik_ELE419_Project__NOR_gate2
Xinverter_1 0 net_30 A_or_B vdd ServetCelik_ELE419_Project__inverter2
.ENDS ServetCelik_ELE419_Project__OR_gate2

*** SUBCIRCUIT ServetCelik_ELE419_Project__NAND_gate2 FROM CELL NAND_gate2{lay}
.SUBCKT ServetCelik_ELE419_Project__NAND_gate2 0 A A_nand_B B vdd
Mnmos_0 net_34 B A_nand_B 0 N L=0.6U W=2.4U AS=4.56P AD=1.418P PS=7.3U PD=4.05U
Mnmos_1 0 A net_34 0 N L=0.6U W=2.4U AS=1.418P AD=16.83P PS=4.05U PD=27.9U
Mpmos_0 A_nand_B A vdd vdd P L=0.6U W=2.4U AS=13.05P AD=4.56P PS=21U PD=7.3U
Mpmos_1 vdd B A_nand_B vdd P L=0.6U W=2.4U AS=4.56P AD=13.05P PS=7.3U PD=21U
.ENDS ServetCelik_ELE419_Project__NAND_gate2

*** SUBCIRCUIT ServetCelik_ELE419_Project__AND_gate2 FROM CELL AND_gate2{lay}
.SUBCKT ServetCelik_ELE419_Project__AND_gate2 0 A A_and_B B vdd
XNAND_gat_2 0 A net_0 B vdd ServetCelik_ELE419_Project__NAND_gate2
Xinverter_2 0 net_0 A_and_B vdd ServetCelik_ELE419_Project__inverter2
.ENDS ServetCelik_ELE419_Project__AND_gate2

*** SUBCIRCUIT ServetCelik_ELE419_Project__XOR_gate2 FROM CELL XOR_gate2{lay}
.SUBCKT ServetCelik_ELE419_Project__XOR_gate2 0 A A_xor_B B vdd
Mnmos_7 net_258 B 0 0 N L=0.6U W=1.2U AS=5.783P AD=1.845P PS=11.7U PD=4.2U
Mnmos_8 A_xor_B A net_258 0 N L=0.6U W=1.2U AS=1.845P AD=2.858P PS=4.2U PD=5.1U
Mnmos_9 net_259 net_263 A_xor_B 0 N L=0.6U W=1.2U AS=2.858P AD=2.025P PS=5.1U PD=4.5U
Mnmos_10 0 net_230 net_259 0 N L=0.6U W=1.2U AS=2.025P AD=5.783P PS=4.5U PD=11.7U
Mnmos_11 net_263 A 0 0 N L=0.6U W=1.2U AS=5.783P AD=4.185P PS=11.7U PD=8.4U
Mnmos_12 net_230 B 0 0 N L=0.6U W=1.2U AS=5.783P AD=4.725P PS=11.7U PD=9U
Mpmos_10 A_xor_B B net_199 vdd P L=0.6U W=2.4U AS=4.995P AD=2.858P PS=8.1U PD=5.1U
Mpmos_11 net_199 A A_xor_B vdd P L=0.6U W=2.4U AS=2.858P AD=4.995P PS=5.1U PD=8.1U
Mpmos_12 vdd net_263 net_199 vdd P L=0.6U W=2.4U AS=4.995P AD=7.808P PS=8.1U PD=12.6U
Mpmos_13 net_199 net_230 vdd vdd P L=0.6U W=2.4U AS=7.808P AD=4.995P PS=12.6U PD=8.1U
Mpmos_14 net_263 A vdd vdd P L=0.6U W=2.4U AS=7.808P AD=4.185P PS=12.6U PD=8.4U
Mpmos_15 net_230 B vdd vdd P L=0.6U W=2.4U AS=7.808P AD=4.725P PS=12.6U PD=9U
.ENDS ServetCelik_ELE419_Project__XOR_gate2

*** SUBCIRCUIT ServetCelik_ELE419_Project__halfAdder2 FROM CELL halfAdder2{lay}
.SUBCKT ServetCelik_ELE419_Project__halfAdder2 0 A B halfAdder_carry halfAdder_sum vdd
XAND_gate_2 0 A halfAdder_carry B vdd ServetCelik_ELE419_Project__AND_gate2
XXOR_gate_2 0 A halfAdder_sum B vdd ServetCelik_ELE419_Project__XOR_gate2
.ENDS ServetCelik_ELE419_Project__halfAdder2

*** SUBCIRCUIT ServetCelik_ELE419_Project__fullAdder2 FROM CELL fullAdder2{lay}
.SUBCKT ServetCelik_ELE419_Project__fullAdder2 0 A B Cin fullAdder_carry fullAdder_sum vdd
XOR_gate2_0 0 net_39 fullAdder_carry net_42 vdd ServetCelik_ELE419_Project__OR_gate2
XhalfAdde_2 0 net_47 Cin net_42 fullAdder_sum vdd ServetCelik_ELE419_Project__halfAdder2
XhalfAdde_3 0 A B net_39 net_47 vdd ServetCelik_ELE419_Project__halfAdder2
.ENDS ServetCelik_ELE419_Project__fullAdder2

*** SUBCIRCUIT ServetCelik_ELE419_Project__2bit_RCA2 FROM CELL 2bit_RCA2{lay}
.SUBCKT ServetCelik_ELE419_Project__2bit_RCA2 0 A0 A1 B0 B1 carry S0 S1 vdd
XfullAdde_2 0 A1 B1 net_34 carry S1 vdd ServetCelik_ELE419_Project__fullAdder2
XfullAdde_3 0 A0 B0 0 net_34 S0 vdd ServetCelik_ELE419_Project__fullAdder2
.ENDS ServetCelik_ELE419_Project__2bit_RCA2

*** SUBCIRCUIT ServetCelik_ELE419_Project__2bit_multiplier2 FROM CELL 2bit_multiplier2{lay}
.SUBCKT ServetCelik_ELE419_Project__2bit_multiplier2 0 A0 A1 B0 B1 P0 P1 P2 P3 vdd
XAND_gate_4 0 A1 net_18 B1 vdd ServetCelik_ELE419_Project__AND_gate2
XAND_gate_5 0 A0 net_11 B1 vdd ServetCelik_ELE419_Project__AND_gate2
XAND_gate_6 0 A1 net_0 B0 vdd ServetCelik_ELE419_Project__AND_gate2
XAND_gate_7 0 A0 P0 B0 vdd ServetCelik_ELE419_Project__AND_gate2
XhalfAdde_2 0 net_11 net_0 net_21 P1 vdd ServetCelik_ELE419_Project__halfAdder2
XhalfAdde_3 0 net_18 net_21 P3 P2 vdd ServetCelik_ELE419_Project__halfAdder2
.ENDS ServetCelik_ELE419_Project__2bit_multiplier2

*** SUBCIRCUIT ServetCelik_ELE419_Project__4bit_RCA2 FROM CELL 4bit_RCA2{lay}
.SUBCKT ServetCelik_ELE419_Project__4bit_RCA2 0 A0 A1 A2 A3 B0 B1 B2 B3 carry S0 S1 S2 S3 vdd
XfullAdde_4 0 A1 B1 net_175 net_106 S1 vdd ServetCelik_ELE419_Project__fullAdder2
XfullAdde_5 0 A0 B0 0 net_175 S0 vdd ServetCelik_ELE419_Project__fullAdder2
XfullAdde_8 0 A3 B3 net_208 carry S3 vdd ServetCelik_ELE419_Project__fullAdder2
XfullAdde_9 0 A2 B2 net_106 net_208 S2 vdd ServetCelik_ELE419_Project__fullAdder2
.ENDS ServetCelik_ELE419_Project__4bit_RCA2

*** SUBCIRCUIT ServetCelik_ELE419_Project__4bit_multiplier2 FROM CELL 4bit_multiplier2{lay}
.SUBCKT ServetCelik_ELE419_Project__4bit_multiplier2 0 A0 A1 A2 A3 B0 B1 B2 B3 carry P0 P1 P2 P3 P4 P5 P6 P7 vdd
X2bit_RCA_1 0 net_762 net_755 net_771 net_783 carry P6 P7 vdd ServetCelik_ELE419_Project__2bit_RCA2
X2bit_mul_4 0 A2 A3 B2 B3 net_369 net_364 net_771 net_783 vdd ServetCelik_ELE419_Project__2bit_multiplier2
X2bit_mul_5 0 A0 A1 B2 B3 net_249 net_258 net_311 net_316 vdd ServetCelik_ELE419_Project__2bit_multiplier2
X2bit_mul_6 0 A2 A3 B0 B1 net_288 net_291 net_296 net_299 vdd ServetCelik_ELE419_Project__2bit_multiplier2
X2bit_mul_7 0 A0 A1 B0 B1 P0 P1 net_350 net_353 vdd ServetCelik_ELE419_Project__2bit_multiplier2
X4bit_RCA_2 0 net_288 net_291 net_296 net_299 net_249 net_258 net_311 net_316 net_752 net_322 net_326 net_330 net_335 vdd ServetCelik_ELE419_Project__4bit_RCA2
X4bit_RCA_3 0 net_350 net_353 net_369 net_364 net_322 net_326 net_330 net_335 net_743 P2 P3 P4 P5 vdd ServetCelik_ELE419_Project__4bit_RCA2
XhalfAdde_2 0 net_752 net_743 net_755 net_762 vdd ServetCelik_ELE419_Project__halfAdder2
.ENDS ServetCelik_ELE419_Project__4bit_multiplier2

*** SUBCIRCUIT ServetCelik_ELE419_Project__3in_NAND_gate2 FROM CELL 3in_NAND_gate2{lay}
.SUBCKT ServetCelik_ELE419_Project__3in_NAND_gate2 0 A A_B_C_nand B C vdd
Mnmos_0 net_34 B net_55 0 N L=0.6U W=3.6U AS=1.958P AD=1.958P PS=5.25U PD=5.25U
Mnmos_1 0 A net_34 0 N L=0.6U W=3.6U AS=1.958P AD=19.62P PS=5.25U PD=30.9U
Mnmos_2 net_55 C A_B_C_nand 0 N L=0.6U W=3.6U AS=5.962P AD=1.958P PS=9U PD=5.25U
Mpmos_0 A_B_C_nand A vdd vdd P L=0.6U W=2.4U AS=9.06P AD=5.962P PS=14.3U PD=9U
Mpmos_1 vdd B A_B_C_nand vdd P L=0.6U W=2.4U AS=5.962P AD=9.06P PS=9U PD=14.3U
Mpmos_2 A_B_C_nand C vdd vdd P L=0.6U W=2.4U AS=9.06P AD=5.962P PS=14.3U PD=9U
.ENDS ServetCelik_ELE419_Project__3in_NAND_gate2

*** SUBCIRCUIT ServetCelik_ELE419_Project__3in_and FROM CELL 3in_and{lay}
.SUBCKT ServetCelik_ELE419_Project__3in_and 0 A ABC_and B C vdd
X3in_NAND_0 0 C net_16 B A vdd ServetCelik_ELE419_Project__3in_NAND_gate2
Xinverter_0 0 net_16 ABC_and vdd ServetCelik_ELE419_Project__inverter2
.ENDS ServetCelik_ELE419_Project__3in_and

*** SUBCIRCUIT ServetCelik_ELE419_Project__8bit_ADD_SUB FROM CELL 8bit_ADD_SUB{lay}
.SUBCKT ServetCelik_ELE419_Project__8bit_ADD_SUB 0 A0 A1 A2 A3 A4 A5 A6 A7 B0 B1 B2 B3 B4 B5 B6 B7 carry Op0 Op1 Op2 S0 S1 S2 S3 S4 S5 S6 S7 vdd
X3in_and_0 0 Op0 net_380 Op1 Op2 vdd ServetCelik_ELE419_Project__3in_and
XXOR_gate_0 0 net_380 net_406 B0 vdd ServetCelik_ELE419_Project__XOR_gate2
XXOR_gate_1 0 net_380 net_142 B1 vdd ServetCelik_ELE419_Project__XOR_gate2
XXOR_gate_2 0 net_380 net_193 B4 vdd ServetCelik_ELE419_Project__XOR_gate2
XXOR_gate_3 0 net_380 net_131 B2 vdd ServetCelik_ELE419_Project__XOR_gate2
XXOR_gate_4 0 net_380 net_201 B6 vdd ServetCelik_ELE419_Project__XOR_gate2
XXOR_gate_5 0 net_380 net_212 B5 vdd ServetCelik_ELE419_Project__XOR_gate2
XXOR_gate_6 0 net_380 net_133 B3 vdd ServetCelik_ELE419_Project__XOR_gate2
XXOR_gate_7 0 net_380 net_203 B7 vdd ServetCelik_ELE419_Project__XOR_gate2
XfullAdde_8 0 A1 net_142 net_139 net_126 S1 vdd ServetCelik_ELE419_Project__fullAdder2
XfullAdde_9 0 A0 net_406 net_380 net_139 S0 vdd ServetCelik_ELE419_Project__fullAdder2
XfullAdde_10 0 A3 net_133 net_165 net_263 S3 vdd ServetCelik_ELE419_Project__fullAdder2
XfullAdde_11 0 A2 net_131 net_126 net_165 S2 vdd ServetCelik_ELE419_Project__fullAdder2
XfullAdde_12 0 A5 net_212 net_209 net_196 S5 vdd ServetCelik_ELE419_Project__fullAdder2
XfullAdde_13 0 A4 net_193 net_263 net_209 S4 vdd ServetCelik_ELE419_Project__fullAdder2
XfullAdde_14 0 A7 net_203 net_235 carry S7 vdd ServetCelik_ELE419_Project__fullAdder2
XfullAdde_15 0 A6 net_201 net_196 net_235 S6 vdd ServetCelik_ELE419_Project__fullAdder2
.ENDS ServetCelik_ELE419_Project__8bit_ADD_SUB

*** SUBCIRCUIT ServetCelik_ELE419_Project__2x1MUX_2 FROM CELL 2x1MUX_2{lay}
.SUBCKT ServetCelik_ELE419_Project__2x1MUX_2 0 D0 D1 OpCode0 out vdd
XAND_gate_0 0 net_106 net_146 D0 vdd ServetCelik_ELE419_Project__AND_gate2
XAND_gate_1 0 OpCode0 net_143 D1 vdd ServetCelik_ELE419_Project__AND_gate2
XOR_gate2_0 0 net_143 out net_146 vdd ServetCelik_ELE419_Project__OR_gate2
Xinverter_0 0 OpCode0 net_106 vdd ServetCelik_ELE419_Project__inverter2
.ENDS ServetCelik_ELE419_Project__2x1MUX_2

*** SUBCIRCUIT ServetCelik_ELE419_Project__8bit_Shifter FROM CELL 8bit_Shifter{lay}
.SUBCKT ServetCelik_ELE419_Project__8bit_Shifter 0 D0 D1 D2 D3 D4 D5 D6 D7 Op0 Op1 S0 S1 S2 S3 S4 S5 S6 S7 vdd
X2x1MUX_2_0 0 net_67 net_72 Op0 S7 vdd ServetCelik_ELE419_Project__2x1MUX_2
X2x1MUX_2_1 0 net_62 net_67 Op0 S6 vdd ServetCelik_ELE419_Project__2x1MUX_2
X2x1MUX_2_2 0 net_57 net_62 Op0 S5 vdd ServetCelik_ELE419_Project__2x1MUX_2
X2x1MUX_2_3 0 net_52 net_57 Op0 S4 vdd ServetCelik_ELE419_Project__2x1MUX_2
X2x1MUX_2_4 0 net_47 net_52 Op0 S3 vdd ServetCelik_ELE419_Project__2x1MUX_2
X2x1MUX_2_5 0 net_41 net_47 Op0 S2 vdd ServetCelik_ELE419_Project__2x1MUX_2
X2x1MUX_2_6 0 net_35 net_41 Op0 S1 vdd ServetCelik_ELE419_Project__2x1MUX_2
X2x1MUX_2_7 0 net_143 net_35 Op0 S0 vdd ServetCelik_ELE419_Project__2x1MUX_2
X2x1MUX_2_8 0 D7 0 Op1 net_72 vdd ServetCelik_ELE419_Project__2x1MUX_2
X2x1MUX_2_9 0 D6 0 Op1 net_67 vdd ServetCelik_ELE419_Project__2x1MUX_2
X2x1MUX_2_10 0 D5 D7 Op1 net_62 vdd ServetCelik_ELE419_Project__2x1MUX_2
X2x1MUX_2_11 0 D4 D6 Op1 net_57 vdd ServetCelik_ELE419_Project__2x1MUX_2
X2x1MUX_2_12 0 D3 D5 Op1 net_52 vdd ServetCelik_ELE419_Project__2x1MUX_2
X2x1MUX_2_13 0 D2 D4 Op1 net_47 vdd ServetCelik_ELE419_Project__2x1MUX_2
X2x1MUX_2_14 0 D1 D3 Op1 net_41 vdd ServetCelik_ELE419_Project__2x1MUX_2
X2x1MUX_2_15 0 D0 D2 Op1 net_35 vdd ServetCelik_ELE419_Project__2x1MUX_2
X2x1MUX_2_16 0 0 D1 Op1 net_143 vdd ServetCelik_ELE419_Project__2x1MUX_2
.ENDS ServetCelik_ELE419_Project__8bit_Shifter

*** SUBCIRCUIT ServetCelik_ELE419_Project__2x1MUX FROM CELL 2x1MUX{lay}
.SUBCKT ServetCelik_ELE419_Project__2x1MUX 0 D0 D1 OpCode0 out vdd
XAND_gate_0 0 net_106 net_146 D0 vdd ServetCelik_ELE419_Project__AND_gate2
XAND_gate_1 0 OpCode0 net_143 D1 vdd ServetCelik_ELE419_Project__AND_gate2
XOR_gate2_0 0 net_143 out net_146 vdd ServetCelik_ELE419_Project__OR_gate2
Xinverter_0 0 OpCode0 net_106 vdd ServetCelik_ELE419_Project__inverter2
.ENDS ServetCelik_ELE419_Project__2x1MUX

*** SUBCIRCUIT ServetCelik_ELE419_Project__4x1MUX FROM CELL 4x1MUX{lay}
.SUBCKT ServetCelik_ELE419_Project__4x1MUX 0 4x1MUX_out D0 D1 D2 D3 OpCode0 OpCode1 vdd
X3in_and_0 0 net_18 net_70 net_3 D0 vdd ServetCelik_ELE419_Project__3in_and
X3in_and_1 0 OpCode0 net_67 net_18 D1 vdd ServetCelik_ELE419_Project__3in_and
X3in_and_2 0 OpCode1 net_77 net_3 D2 vdd ServetCelik_ELE419_Project__3in_and
X3in_and_3 0 OpCode0 net_74 OpCode1 D3 vdd ServetCelik_ELE419_Project__3in_and
XOR_gate2_0 0 net_67 net_81 net_70 vdd ServetCelik_ELE419_Project__OR_gate2
XOR_gate2_1 0 net_74 net_85 net_77 vdd ServetCelik_ELE419_Project__OR_gate2
XOR_gate2_2 0 net_85 4x1MUX_out net_81 vdd ServetCelik_ELE419_Project__OR_gate2
Xinverter_0 0 OpCode0 net_3 vdd ServetCelik_ELE419_Project__inverter2
Xinverter_1 0 OpCode1 net_18 vdd ServetCelik_ELE419_Project__inverter2
.ENDS ServetCelik_ELE419_Project__4x1MUX

*** SUBCIRCUIT ServetCelik_ELE419_Project__8x1MUX FROM CELL 8x1MUX{lay}
.SUBCKT ServetCelik_ELE419_Project__8x1MUX 0 D0 D1 D2 D3 D4 D5 D6 D7 OpCode0 OpCode1 OpCode2 Out vdd
X2x1MUX_0 0 net_91 net_89 OpCode2 Out vdd ServetCelik_ELE419_Project__2x1MUX
X4x1MUX_0 0 net_91 D0 D1 D2 D3 OpCode0 OpCode1 vdd ServetCelik_ELE419_Project__4x1MUX
X4x1MUX_1 0 net_89 D4 D5 D6 D7 OpCode0 OpCode1 vdd ServetCelik_ELE419_Project__4x1MUX
.ENDS ServetCelik_ELE419_Project__8x1MUX

*** SUBCIRCUIT ServetCelik_ELE419_Project__8x1MUX_8bit FROM CELL 8x1MUX_8bit{lay}
.SUBCKT ServetCelik_ELE419_Project__8x1MUX_8bit 0 B00 B01 B02 B03 B04 B05 B06 B07 B10 B11 B12 B13 B14 B15 B16 B17 B20 B21 B22 B23 B24 B25 B26 B27 B31 B32 B33 B34 B35 B36 B37 B40 B41 B42 B43 B44 B45 B46 B47 B50 B51 B52 B53 B54 B55 B56 B57 B60 B61 B62 B63 B64 B65 B66 B67 B70 B71 B72 B73 B74 B75 B76 B77 OpCode0 OpCode1 OpCode2 Out0 Out1 Out2 Out3 Out4 Out5 Out6 Out7 V30 vdd
X8x1MUX_0 0 B70 B71 B72 B73 B74 B75 B76 B77 OpCode0 OpCode1 OpCode2 Out7 vdd ServetCelik_ELE419_Project__8x1MUX
X8x1MUX_1 0 B60 B61 B62 B63 B64 B65 B66 B67 OpCode0 OpCode1 OpCode2 Out6 vdd ServetCelik_ELE419_Project__8x1MUX
X8x1MUX_2 0 B50 B51 B52 B53 B54 B55 B56 B57 OpCode0 OpCode1 OpCode2 Out5 vdd ServetCelik_ELE419_Project__8x1MUX
X8x1MUX_3 0 B40 B41 B42 B43 B44 B45 B46 B47 OpCode0 OpCode1 OpCode2 Out4 vdd ServetCelik_ELE419_Project__8x1MUX
X8x1MUX_4 0 V30 B31 B32 B33 B34 B35 B36 B37 OpCode0 OpCode1 OpCode2 Out3 vdd ServetCelik_ELE419_Project__8x1MUX
X8x1MUX_5 0 B20 B21 B22 B23 B24 B25 B26 B27 OpCode0 OpCode1 OpCode2 Out2 vdd ServetCelik_ELE419_Project__8x1MUX
X8x1MUX_6 0 B10 B11 B12 B13 B14 B15 B16 B17 OpCode0 OpCode1 OpCode2 Out1 vdd ServetCelik_ELE419_Project__8x1MUX
X8x1MUX_7 0 B00 B01 B02 B03 B04 B05 B06 B07 OpCode0 OpCode1 OpCode2 Out0 vdd ServetCelik_ELE419_Project__8x1MUX
.ENDS ServetCelik_ELE419_Project__8x1MUX_8bit

*** SUBCIRCUIT ServetCelik_ELE419_Project__inverter_8bit FROM CELL inverter_8bit{lay}
.SUBCKT ServetCelik_ELE419_Project__inverter_8bit 0 A0 A1 A2 A3 A4 A5 A6 A7 S0 S1 S2 S3 S4 S5 S6 S7 vdd
Xinverter_0 0 A7 S7 vdd ServetCelik_ELE419_Project__inverter2
Xinverter_1 0 A6 S6 vdd ServetCelik_ELE419_Project__inverter2
Xinverter_2 0 A5 S5 vdd ServetCelik_ELE419_Project__inverter2
Xinverter_3 0 A4 S4 vdd ServetCelik_ELE419_Project__inverter2
Xinverter_8 0 A3 S3 vdd ServetCelik_ELE419_Project__inverter2
Xinverter_9 0 A2 S2 vdd ServetCelik_ELE419_Project__inverter2
Xinverter_10 0 A1 S1 vdd ServetCelik_ELE419_Project__inverter2
Xinverter_11 0 A0 S0 vdd ServetCelik_ELE419_Project__inverter2
.ENDS ServetCelik_ELE419_Project__inverter_8bit

*** TOP LEVEL CELL: 8bit_ALU{lay}
X4bit_mul_0 0 A0 A1 A2 A3 B0 B1 B2 B3 4bit_mul_0_carry net_570 net_573 net_576 net_579 net_582 net_585 net_588 net_591 vdd ServetCelik_ELE419_Project__4bit_multiplier2
X8bit_ADD_0 0 A0 A1 A2 A3 A4 A5 A6 A7 B0 B1 B2 B3 B4 B5 B6 B7 8bit_ADD_0_carry OpCode0 OpCode1 OpCode2 net_281 net_284 net_287 net_290 net_292 net_295 net_298 net_301 vdd ServetCelik_ELE419_Project__8bit_ADD_SUB
X8bit_Shi_0 0 A0 A1 A2 A3 A4 A5 A6 A7 OpCode0 OpCode1 net_130 net_136 net_139 net_142 net_145 net_148 net_151 net_154 vdd ServetCelik_ELE419_Project__8bit_Shifter
X8x1MUX_8_0 0 net_130 net_130 net_130 net_130 net_570 net_537 net_281 net_281 net_136 net_136 net_136 net_136 net_573 net_639 net_284 net_284 net_139 net_139 net_139 net_139 net_576 net_636 net_287 net_287 net_142 net_142 net_142 net_579 net_633 net_290 net_290 net_145 net_145 net_145 net_145 net_582 net_629 net_292 net_292 net_148 net_148 net_148 net_148 net_585 net_626 net_295 net_295 net_151 net_151 net_151 net_151 net_588 net_623 net_298 net_298 net_154 net_154 net_154 net_154 net_591 net_621 net_301 
+net_301 OpCode0 OpCode1 OpCode2 Out0 Out1 Out2 Out3 Out4 Out5 Out6 Out7 net_142 vdd ServetCelik_ELE419_Project__8x1MUX_8bit
Xinverter_0 0 A0 A1 A2 A3 A4 A5 A6 A7 net_537 net_639 net_636 net_633 net_629 net_626 net_623 net_621 vdd ServetCelik_ELE419_Project__inverter_8bit

* Spice Code nodes in cell cell '8bit_ALU{lay}'
vdd vdd 0 DC 5
VinOpCode0 OpCode0 0 DC 0
VinOpCode1 OpCode1 0 DC 0
VinOpCode2 OpCode2 0 DC 0
VinA7 A7 0 DC 5
VinA6 A6 0 DC 0
VinA5 A5 0 DC 0
VinA4 A4 0 DC 5
VinA3 A3 0 DC 0
VinA2 A2 0 DC 0
VinA1 A1 0 DC 0
VinA0 A0 0 DC 5
.tran 10u 40u
* Trailer cards are described in this file:
.INC C:\Users\Servet\Desktop\C5_models.txt
.END
