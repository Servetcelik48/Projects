*** SPICE deck for cell 8bit_ADD_SUB{lay} from library ServetCelik_ELE419_Project
*** Created on Pzt Oca 01, 2024 22:50:46
*** Last revised on Pzt Oca 15, 2024 08:31:10
*** Written on Pzt Oca 15, 2024 08:31:17 by Electric VLSI Design System, version 9.07
*** Layout tech: mocmos, foundry MOSIS
*** UC SPICE *** , MIN_RESIST 4.0, MIN_CAPAC 0.1FF

*** SUBCIRCUIT ServetCelik_ELE419_Project__3in_NAND_gate2 FROM CELL 3in_NAND_gate2{lay}
.SUBCKT ServetCelik_ELE419_Project__3in_NAND_gate2 0 A A_B_C_nand B C vdd
Mnmos_0 net_34 B net_55 0 N L=0.6U W=3.6U AS=1.958P AD=1.958P PS=5.25U PD=5.25U
Mnmos_1 0 A net_34 0 N L=0.6U W=3.6U AS=1.958P AD=19.62P PS=5.25U PD=30.9U
Mnmos_2 net_55 C A_B_C_nand 0 N L=0.6U W=3.6U AS=5.962P AD=1.958P PS=9U PD=5.25U
Mpmos_0 A_B_C_nand A vdd vdd P L=0.6U W=2.4U AS=9.06P AD=5.962P PS=14.3U PD=9U
Mpmos_1 vdd B A_B_C_nand vdd P L=0.6U W=2.4U AS=5.962P AD=9.06P PS=9U PD=14.3U
Mpmos_2 A_B_C_nand C vdd vdd P L=0.6U W=2.4U AS=9.06P AD=5.962P PS=14.3U PD=9U
.ENDS ServetCelik_ELE419_Project__3in_NAND_gate2

*** SUBCIRCUIT ServetCelik_ELE419_Project__inverter2 FROM CELL inverter2{lay}
.SUBCKT ServetCelik_ELE419_Project__inverter2 0 A A_not vdd
Mnmos_0 A_not A 0 0 N L=0.6U W=1.2U AS=9.54P AD=4.725P PS=18.9U PD=9U
Mpmos_0 A_not A vdd vdd P L=0.6U W=2.4U AS=12.33P AD=4.725P PS=21.9U PD=9U
.ENDS ServetCelik_ELE419_Project__inverter2

*** SUBCIRCUIT ServetCelik_ELE419_Project__3in_and FROM CELL 3in_and{lay}
.SUBCKT ServetCelik_ELE419_Project__3in_and 0 A ABC_and B C vdd
X3in_NAND_0 0 C net_16 B A vdd ServetCelik_ELE419_Project__3in_NAND_gate2
Xinverter_0 0 net_16 ABC_and vdd ServetCelik_ELE419_Project__inverter2
.ENDS ServetCelik_ELE419_Project__3in_and

*** SUBCIRCUIT ServetCelik_ELE419_Project__XOR_gate2 FROM CELL XOR_gate2{lay}
.SUBCKT ServetCelik_ELE419_Project__XOR_gate2 0 A A_xor_B B vdd
Mnmos_7 net_258 B 0 0 N L=0.6U W=1.2U AS=5.783P AD=1.845P PS=11.7U PD=4.2U
Mnmos_8 A_xor_B A net_258 0 N L=0.6U W=1.2U AS=1.845P AD=2.858P PS=4.2U PD=5.1U
Mnmos_9 net_259 net_263 A_xor_B 0 N L=0.6U W=1.2U AS=2.858P AD=2.025P PS=5.1U PD=4.5U
Mnmos_10 0 net_230 net_259 0 N L=0.6U W=1.2U AS=2.025P AD=5.783P PS=4.5U PD=11.7U
Mnmos_11 net_263 A 0 0 N L=0.6U W=1.2U AS=5.783P AD=4.185P PS=11.7U PD=8.4U
Mnmos_12 net_230 B 0 0 N L=0.6U W=1.2U AS=5.783P AD=4.725P PS=11.7U PD=9U
Mpmos_10 A_xor_B B net_199 vdd P L=0.6U W=2.4U AS=4.995P AD=2.858P PS=8.1U PD=5.1U
Mpmos_11 net_199 A A_xor_B vdd P L=0.6U W=2.4U AS=2.858P AD=4.995P PS=5.1U PD=8.1U
Mpmos_12 vdd net_263 net_199 vdd P L=0.6U W=2.4U AS=4.995P AD=7.808P PS=8.1U PD=12.6U
Mpmos_13 net_199 net_230 vdd vdd P L=0.6U W=2.4U AS=7.808P AD=4.995P PS=12.6U PD=8.1U
Mpmos_14 net_263 A vdd vdd P L=0.6U W=2.4U AS=7.808P AD=4.185P PS=12.6U PD=8.4U
Mpmos_15 net_230 B vdd vdd P L=0.6U W=2.4U AS=7.808P AD=4.725P PS=12.6U PD=9U
.ENDS ServetCelik_ELE419_Project__XOR_gate2

*** SUBCIRCUIT ServetCelik_ELE419_Project__NOR_gate2 FROM CELL NOR_gate2{lay}
.SUBCKT ServetCelik_ELE419_Project__NOR_gate2 0 A A_nor_B B vdd
Mnmos_2 A_nor_B A 0 0 N L=0.6U W=1.2U AS=6.525P AD=3.21P PS=13.5U PD=6.1U
Mnmos_3 0 B A_nor_B 0 N L=0.6U W=1.2U AS=3.21P AD=6.525P PS=6.1U PD=13.5U
Mpmos_2 net_75 A vdd vdd P L=0.6U W=2.4U AS=13.05P AD=1.418P PS=22.5U PD=4.05U
Mpmos_3 A_nor_B B net_75 vdd P L=0.6U W=2.4U AS=1.418P AD=3.21P PS=4.05U PD=6.1U
.ENDS ServetCelik_ELE419_Project__NOR_gate2

*** SUBCIRCUIT ServetCelik_ELE419_Project__OR_gate2 FROM CELL OR_gate2{lay}
.SUBCKT ServetCelik_ELE419_Project__OR_gate2 0 A A_or_B B vdd
XNOR_gate_2 0 A net_30 B vdd ServetCelik_ELE419_Project__NOR_gate2
Xinverter_1 0 net_30 A_or_B vdd ServetCelik_ELE419_Project__inverter2
.ENDS ServetCelik_ELE419_Project__OR_gate2

*** SUBCIRCUIT ServetCelik_ELE419_Project__NAND_gate2 FROM CELL NAND_gate2{lay}
.SUBCKT ServetCelik_ELE419_Project__NAND_gate2 0 A A_nand_B B vdd
Mnmos_0 net_34 B A_nand_B 0 N L=0.6U W=2.4U AS=4.56P AD=1.418P PS=7.3U PD=4.05U
Mnmos_1 0 A net_34 0 N L=0.6U W=2.4U AS=1.418P AD=16.83P PS=4.05U PD=27.9U
Mpmos_0 A_nand_B A vdd vdd P L=0.6U W=2.4U AS=13.05P AD=4.56P PS=21U PD=7.3U
Mpmos_1 vdd B A_nand_B vdd P L=0.6U W=2.4U AS=4.56P AD=13.05P PS=7.3U PD=21U
.ENDS ServetCelik_ELE419_Project__NAND_gate2

*** SUBCIRCUIT ServetCelik_ELE419_Project__AND_gate2 FROM CELL AND_gate2{lay}
.SUBCKT ServetCelik_ELE419_Project__AND_gate2 0 A A_and_B B vdd
XNAND_gat_2 0 A net_0 B vdd ServetCelik_ELE419_Project__NAND_gate2
Xinverter_2 0 net_0 A_and_B vdd ServetCelik_ELE419_Project__inverter2
.ENDS ServetCelik_ELE419_Project__AND_gate2

*** SUBCIRCUIT ServetCelik_ELE419_Project__halfAdder2 FROM CELL halfAdder2{lay}
.SUBCKT ServetCelik_ELE419_Project__halfAdder2 0 A B halfAdder_carry halfAdder_sum vdd
XAND_gate_2 0 A halfAdder_carry B vdd ServetCelik_ELE419_Project__AND_gate2
XXOR_gate_2 0 A halfAdder_sum B vdd ServetCelik_ELE419_Project__XOR_gate2
.ENDS ServetCelik_ELE419_Project__halfAdder2

*** SUBCIRCUIT ServetCelik_ELE419_Project__fullAdder2 FROM CELL fullAdder2{lay}
.SUBCKT ServetCelik_ELE419_Project__fullAdder2 0 A B Cin fullAdder_carry fullAdder_sum vdd
XOR_gate2_0 0 net_39 fullAdder_carry net_42 vdd ServetCelik_ELE419_Project__OR_gate2
XhalfAdde_2 0 net_47 Cin net_42 fullAdder_sum vdd ServetCelik_ELE419_Project__halfAdder2
XhalfAdde_3 0 A B net_39 net_47 vdd ServetCelik_ELE419_Project__halfAdder2
.ENDS ServetCelik_ELE419_Project__fullAdder2

*** TOP LEVEL CELL: 8bit_ADD_SUB{lay}
X3in_and_0 0 vdd net_380 vdd vdd vdd ServetCelik_ELE419_Project__3in_and
XXOR_gate_0 0 net_380 net_406 B0 vdd ServetCelik_ELE419_Project__XOR_gate2
XXOR_gate_1 0 net_380 net_142 B1 vdd ServetCelik_ELE419_Project__XOR_gate2
XXOR_gate_2 0 net_380 net_193 B4 vdd ServetCelik_ELE419_Project__XOR_gate2
XXOR_gate_3 0 net_380 net_131 B2 vdd ServetCelik_ELE419_Project__XOR_gate2
XXOR_gate_4 0 net_380 net_201 B6 vdd ServetCelik_ELE419_Project__XOR_gate2
XXOR_gate_5 0 net_380 net_212 B5 vdd ServetCelik_ELE419_Project__XOR_gate2
XXOR_gate_6 0 net_380 net_133 B3 vdd ServetCelik_ELE419_Project__XOR_gate2
XXOR_gate_7 0 net_380 net_203 B7 vdd ServetCelik_ELE419_Project__XOR_gate2
XfullAdde_8 0 A1 net_142 net_139 net_126 S1 vdd ServetCelik_ELE419_Project__fullAdder2
XfullAdde_9 0 A0 net_406 vdd net_139 S0 vdd ServetCelik_ELE419_Project__fullAdder2
XfullAdde_10 0 A3 net_133 net_165 net_263 S3 vdd ServetCelik_ELE419_Project__fullAdder2
XfullAdde_11 0 A2 net_131 net_126 net_165 S2 vdd ServetCelik_ELE419_Project__fullAdder2
XfullAdde_12 0 A5 net_212 net_209 net_196 S5 vdd ServetCelik_ELE419_Project__fullAdder2
XfullAdde_13 0 A4 net_193 net_263 net_209 S4 vdd ServetCelik_ELE419_Project__fullAdder2
XfullAdde_14 0 A7 net_203 net_235 carry S7 vdd ServetCelik_ELE419_Project__fullAdder2
XfullAdde_15 0 A6 net_201 net_196 net_235 S6 vdd ServetCelik_ELE419_Project__fullAdder2

* Spice Code nodes in cell cell '8bit_ADD_SUB{lay}'
vdd vdd 0 DC 5
VinA7 A7 0 DC 0
VinA6 A6 0 DC 0
VinA5 A5 0 DC 0
VinA4 A4 0 DC 0
VinA3 A3 0 DC 5
VinA2 A2 0 DC 5
VinA1 A1 0 DC 5
VinA0 A0 0 DC 5
VinB7 B7 0 DC 5
VinB6 B6 0 DC 0
VinB5 B5 0 DC 5
VinB4 B4 0 DC 0
VinB3 B3 0 DC 5
VinB2 B2 0 DC 0
VinB1 B1 0 DC 5
VinB0 B0 0 DC 0
.tran 10u 40u
* Trailer cards are described in this file:
.INC C:\Users\Servet\Desktop\C5_models.txt
.END
